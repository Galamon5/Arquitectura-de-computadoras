LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;
LIBRARY MACHXO2;
USE MACHXO2.ALL;

PACKAGE packagemult4bit00 IS
	COMPONENT topfa00
		PORT(C00, B00, A00 : IN STD_LOGIC;
			 S00, C01 : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT and00
		PORT(Aa, Ba : IN STD_LOGIC;
			 Ya     : OUT STD_LOGIC
		 );
	END COMPONENT;
END packagemult4bit00;